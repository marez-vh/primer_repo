library ieee;
use ieee.std_logic_1164.all;
entity example1 is
port(x1, x2 : in std_logic_vector(3 downto 0);
displays: out std_logic_vector(13 downto 0) );
end example1;
architecture bev of example1
begin
--TODO
end bev;